library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;

entity OR_16 is
   port(x_or,y_or: in std_logic_vector(15 downto 0);
	
	s0_or: out std_logic_vector(15 downto 0));
end entity;

architecture Struct of OR_16 is

begin
s0_or<= (x_or or y_or);
end Struct;